`ifndef _RAMmemoryparam_vh_
`define _RAMmemoryparam_vh_
`define RAM_ADDR_BITS 16
`endif