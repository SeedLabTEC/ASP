`ifndef _ROMmemoryparam_vh 
`define _ROMmemoryparam_vh 
`define ROM_ADDR_BITS 12
`define ROM_ADDR_START_BITS 15
`define BEGIN_ADDR_ROM_PROGRAM 32'd32768
`define END_ADDR_ROM_PROGRAM 32'd36863
`define StackPointer 32'd32768
`define ProgramStartAddressPC 32'd32926
`endif